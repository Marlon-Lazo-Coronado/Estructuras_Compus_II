module tournament #(parameter n=32, size=16)( //El alto de la tabla es (2**size)-1
			input reset,
			input clock,
			input fix_result,
			input [n-1:0]etiqueta,
			input [n-1:0]PC,
			output reg [n-1:0]nex_PC,
			output reg prediction);

reg [1:0]table_states[0:1000];
integer i;
reg [1:0]swich;
reg [n-1:0]miss;
reg [n-1:0]hit;

//Logica combinacional
always @(*) begin

	if (reset) begin
		swich[1:0] = 2'b00;
		miss[n-1:0] = 32'h00000000;
		hit[n-1:0] = 32'h00000000;
		
		for (i=0; i<=(2^size)-1; i++)
			table_states [i] = 2'b00;
	end
	else begin
		swich = table_states[PC];
		if ( swich == 2'b00 || swich == 2'b01)begin 
			nex_PC = PC+32'h00000004;
			prediction = 1'b0;
		end
		else begin
			nex_PC = PC+etiqueta;
			prediction = 1'b1;
		end	
	

		//Actualizar el BHT, planteamos varios casos, esto se hace instantaneo, el despase de tiempo lodebe de traer fix_result
		if (fix_result == 1 && prediction==0)//Fallamos!
			table_states[PC] = table_states[PC]+1'b1; //Nos acercamos a gshare
		else if (fix_result == 1 && prediction == 1) begin
			if (swich==2'b10)
				table_states[PC] = table_states[PC]+1'b1;
			else
				table_states[PC] = table_states[PC];
		end
		else if (fix_result == 0 && prediction == 0) begin
			if (swich==2'b01)
				table_states[PC] = table_states[PC]-1'b1; 
			else
				table_states[PC] = table_states[PC];
		end
		else
			table_states[PC] = table_states[PC]-1'b1;
			
		if (fix_result == prediction)
			hit = hit+1'b1;
		else
			miss = miss+1'b1;
	end 
end

endmodule
